module rf;

logic[7:0] core[16];

endmodule